
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity ripple_adder_16_tb is
--  Port ( );
end ripple_adder_16_tb;

architecture Behavioral of ripple_adder_16_tb is

begin


end Behavioral;
